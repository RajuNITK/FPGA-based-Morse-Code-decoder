
module display_project(
	clk,
	reset,
	display_vga,
	onn,
	end_of_active_frame,
	end_of_frame,divcntr,

	// dac pins
	vga_blank,					//	VGA BLANK
	vga_c_sync,					//	VGA COMPOSITE SYNC
	vga_h_sync,					//	VGA H_SYNC
	vga_v_sync,					//	VGA V_SYNC
	//vga_data_enable,			// VGA DEN
	vga_red,						//	VGA Red[9:0]
	vga_green,	 				//	VGA Green[9:0]
	vga_blue,	   			//	VGA Blue[9:0]
	//vga_color_data	   	//	VGA Color[9:0] for TRDB_LCM
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/

parameter CW								= 7;

/* Number of pixels */
parameter H_ACTIVE 						= 640;
parameter H_FRONT_PORCH					=  16;
parameter H_SYNC							=  96;
parameter H_BACK_PORCH 					=  48;
parameter H_TOTAL 						= 800;

/* Number of lines */
parameter V_ACTIVE 						= 480;
parameter V_FRONT_PORCH					=  10;
parameter V_SYNC							=   2;
parameter V_BACK_PORCH 					=  33;
parameter V_TOTAL							= 525;

parameter PW								= 10;			// Number of bits for pixels
parameter PIXEL_COUNTER_INCREMENT	= 10'h001;

parameter LW								= 10;			// Number of bits for lines
parameter LINE_COUNTER_INCREMENT		= 10'h001;

/******************************************************************************/


parameter [419:0] o_pic = {
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},
};

parameter [419:0] x_pic = {
{30'b000000001110000000001110000000},
{30'b000000000111000000011100000000},
{30'b000000000011100000111000000000},
{30'b000000000001110001110000000000},
{30'b000000000000111011100000000000},
{30'b000000000000011111000000000000},
{30'b000000000000001110000000000000},
{30'b000000000000011111000000000000},
{30'b000000000000111011100000000000},
{30'b000000000001110001110000000000},
{30'b000000000011100000110000000000},
{30'b000000000111000000011100000000},
{30'b000000001110000000001110000000},
{30'b000000000000000000000000000000},
};

parameter [419:0] I_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
};

parameter [419:0] T_pic = {
{30'b000001111111111111111111110000},
{30'b000001111111111111111111110000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111110000000000000},

};
 

parameter [419:0] U_pic = {
{30'b000000000000000000000000000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},

};


parameter [419:0] A_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000000000000000000000000000},


};

parameter [419:0] B_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},

};


parameter [419:0] E_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},


};


parameter [419:0] C_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},


};


parameter [419:0] D_pic = {
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},

};



parameter [419:0] F_pic = {
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000000000000000000000000000},

};


parameter [419:0] G_pic = {
{30'b000000000000000000000000000000},
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000011111111000000},
{30'b000000011110000011111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},

};



parameter [419:0] H_pic = {
{30'b000000000000000000000000000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000000000000000000000000000},


};

parameter [419:0] Y_pic = {
{30'b000000000000000000000000000000},
{30'b000000011110000000001110000000},
{30'b000000001111000000011100000000},
{30'b000000000111000000111000000000},
{30'b000000000011100001110000000000},
{30'b000000000001110011100000000000},
{30'b000000000000110111000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000011110000000000000},
{30'b000000000000000000000000000000},
};




parameter [419:0] Z_pic = {
{30'b000000111111111111111110000000},
{30'b000000111111111111111110000000},
{30'b000000000000000000001110000000},
{30'b000000000000000000111110000000},
{30'b000000000000000011111100000000},
{30'b000000000000001111110000000000},
{30'b000000000000011111000000000000},
{30'b000000000011111000000000000000},
{30'b000000000111100000000000000000},
{30'b000000001111100000000000000000},
{30'b000000011111000000000000000000},
{30'b000000111111000000000000000000},
{30'b000000111111111111111110000000},
{30'b000000111111111111111110000000},


};


parameter [419:0] J_pic = {
{30'b000000000000000000000000000000},
{30'b000000111111111111111111111111},
{30'b000000111111111111111111111111},
{30'b000000000000000000111110000000},
{30'b000000000000000000111110000000},
{30'b000000000000000000111110000000},
{30'b000000000000000000111110000000},
{30'b000000000000000000111110000000},
{30'b000000000000000000111110000000},
{30'b000000111100000000111110000000},
{30'b000000111100000000111110000000},
{30'b000000111111111111111110000000},
{30'b000000111111111111111110000000},

};


parameter [419:0] K_pic = {
{30'b000000011100000000011100000000},
{30'b000000011100000001110000000000},
{30'b000000011100000111000000000000},
{30'b000000011100011100000000000000},
{30'b000000011101110000000000000000},
{30'b000000011111000000000000000000},
{30'b000000011100000000000000000000},
{30'b000000011111000000000000000000},
{30'b000000011101110000000000000000},
{30'b000000011100011100000000000000},
{30'b000000011100000111000000000000},
{30'b000000011100000001110000000000},
{30'b000000011100000000011100000000},
{30'b000000000000000000000000000000},

};
parameter [419:0] L_pic = {
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},


};


parameter [419:0] P_pic = {
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},

};


parameter [419:0] R_pic = {
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011110000000001111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111000000000000000},
{30'b000000011110111110000000000000},
{30'b000000011110011111000000000000},
{30'b000000011110001111100000000000},
{30'b000000011110000111110000000000},
{30'b000000011110000011111000000000},
};


parameter [419:0] S_pic = {
{30'b000000000000000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011110000000000000000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000011111000000},
{30'b000000000000000000011111000000},
{30'b000000000000000000011111000000},
{30'b000000011111111111111111000000},
{30'b000000011111111111111111000000},
{30'b000000000000000000000000000000},

};



parameter [419:0] M_pic = {
{30'b000000000000000000000000000000},
{30'b000111111111111111111111000000},
{30'b000111111111111111111111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000000000000000000000000000000},

};

parameter [419:0] N_pic = {
{30'b000000000000000000000000000000},
{30'b000111111100000000001111000000},
{30'b000111101110000000001111000000},
{30'b000111100111000000001111000000},
{30'b000111100011100000001111000000},
{30'b000111100001110000001111000000},
{30'b000111100000111000001111000000},
{30'b000111100000011100001111000000},
{30'b000111100000001110001111000000},
{30'b000111100000000111001111000000},
{30'b000111100000000011101111000000},
{30'b000111100000000001111111000000},
{30'b000111100000000000111111000000},
{30'b000000000000000000000000000000},

};

parameter [419:0] Q_pic = {

{30'b000000111111111111111110000000},
{30'b000000111111111111111110000000},
{30'b000000111100000000011110000000},
{30'b000000111100000000011110000000},
{30'b000000111100000000011110000000},
{30'b000000111100000000011110000000},
{30'b000000111100000000011110000000},
{30'b000000111100000000011110000000},
{30'b000000111100001110011110000000},
{30'b000000111100000111011110000000},
{30'b000000111111111111111110000000},
{30'b000000111111111111111110000000},
{30'b000000000000000000111111000000},
{30'b000000000000000000001111110000},
};

parameter [419:0] V_pic = {
{30'b000000000000000000000000000000},
{30'b111100000000000000000000111100},
{30'b011110000000000000000001111000},
{30'b001111000000000000000011110000},
{30'b000111000000000000000111100000},
{30'b000011110000000000001111000000},
{30'b000001111000000000011110000000},
{30'b000000011110000000111100000000},
{30'b000000001111000001111000000000},
{30'b000000000111100011110000000000},
{30'b000000000011100111100000000000},
{30'b000000000001111111000000000000},
{30'b000000000000111110000000000000},
{30'b000000000000111100000000000000},
{30'b000000000000011000000000000000},
};

parameter [419:0] W_pic = {
{30'b000000000000000000000000000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111100000111100001111000000},
{30'b000111111111111111111111000000},
{30'b000111111111111111111111000000},
};
/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/

input						clk;
input						reset;
input						[4:0] display_vga;
input						onn;
output reg           divcntr;

output reg				end_of_active_frame;
output reg				end_of_frame; 

output reg				vga_blank;			//	VGA BLANK
output reg				vga_c_sync;			//	VGA COMPOSITE SYNC
output reg				vga_h_sync;			//	VGA H_SYNC
output reg				vga_v_sync;			//	VGA V_SYNC
//output reg				vga_data_enable;	// VGA DEN
output reg	[CW: 0]	vga_red;				//	VGA Red[9:0]
output reg	[CW: 0]	vga_green;			//	VGA Green[9:0]
output reg	[CW: 0]	vga_blue;  	 		//	VGA Blue[9:0]
//output reg	[CW: 0]	vga_color_data;	//	VGA Color[9:0] for TRDB_LCM


/*****************************************************************************
 *Internal Wires and Registers Declarations                 *
 *****************************************************************************/
reg			[PW:1]	pixel_counter;
reg			[LW:1]	line_counter;

reg						early_hsync_pulse;
reg						early_vsync_pulse;
reg						hsync_pulse;
reg						vsync_pulse;
reg						csync_pulse;

reg						hblanking_pulse;
reg						vblanking_pulse;
reg						blanking_pulse;

// State Machine Registers
//integers
reg [10:0] m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,
          m20,m21,m22,m23,m24,m25,m26;
/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/
always @(posedge clk)
begin
if(reset) divcntr=1'b0;
 else
 divcntr = ~divcntr;
 //div_clk = divcntr;
 end
///////////////////////////////////////////////////////////////////////////////

always @ (negedge divcntr)
begin
	if (reset)
	begin
		vga_c_sync			<= 1'b1;
		vga_blank			<= 1'b1;
		vga_h_sync			<= 1'b1;
		vga_v_sync			<= 1'b1;

		vga_red				<= {(CW + 1){1'b0}};
		vga_green			<= {(CW + 1){1'b0}};
		vga_blue				<= {(CW + 1){1'b0}};
	m1=10'd419;m2=10'd419;m3=10'd419;m4=10'd419;m5=10'd419;m6=10'd419;m7=10'd419;m8=10'd419;m9=10'd419;m10=10'd419;
	m11=10'd419;m12=10'd419;m13=10'd419;m14=10'd419;m15=10'd419;m16=10'd419;m17=10'd419;m18=10'd419;m19=10'd419;
	m21=10'd419;m22=10'd419;m23=10'd419;m24=10'd419;m25=10'd419;m26=10'd419;
	end
	
	else
	
	begin
		vga_blank			<= ~blanking_pulse;
		vga_c_sync			<= ~csync_pulse;
		vga_h_sync			<= ~hsync_pulse;
		vga_v_sync			<= ~vsync_pulse;
		//vga_data_enable	<= ~blanking_pulse;

		if (blanking_pulse)
		begin
			vga_red			<= {(CW + 1){1'b0}};
			vga_green		<= {(CW + 1){1'b0}};
			vga_blue			<= {(CW + 1){1'b0}};

		end
	
		else
		begin
		///////////////////////////////////////////Display #
		
				/*if((pixel_counter >= 10'd0 && pixel_counter <= 10'd639)  && (line_counter >= 10'd0 && line_counter <= 10'd479)) 
					begin
						//if((pixel_counter > 10'd0 && pixel_counter <= 10'd60)  && (line_counter > 10'd31 && line_counter <= 10'd79))
						//begin
							vga_red<= 8'd0;
							vga_blue<= 8'd255;
							vga_green<= 8'd0;
							end
						//end	*/
				/*if((pixel_counter >= 10'd211 && pixel_counter <= 10'd215) ||
			          (pixel_counter >= 10'd424 && pixel_counter <= 10'd428) ||
						 (line_counter >= 10'd158 && line_counter <= 10'd162) ||
						 (line_counter >= 10'd318 && line_counter <= 10'd322))			
		begin
			vga_red<= 8'd255;
			vga_blue<= 8'd0;
			vga_green<= 8'd0;
		end*/
		
	if((pixel_counter > 10'd30 && pixel_counter <= 10'd60)  && (line_counter > 10'd20 && line_counter <= 10'd34))
			begin
			if(display_vga==5'b00001)
										begin
											if(B_pic[m2])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m2<=m2-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m2==0)
												m2<=10'd419;
												else
												m2<=m2-1'b1;
												
											end
										end
					else if(display_vga==5'b00000)
										begin
											if(A_pic[m1])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m1<=m1-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m1==0)
												m1<=10'd419;
												else
												m1<=m1-1'b1;
												
											end
											end
												else if(display_vga==5'b00010)
										begin
											if(C_pic[m3])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m3<=m3-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m3==0)
												m3<=10'd419;
												else
												m3<=m3-1'b1;
												
											end
											end
												else if(display_vga==5'b00011)
										begin
											if(D_pic[m4])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m4<=m4-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m4==0)
												m4<=10'd419;
												else
												m4<=m4-1'b1;
												
											end
											end
												else if(display_vga==5'b00101)
										begin
											if(E_pic[m5])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m5<=m5-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m5==0)
												m1<=10'd419;
												else
												m5<=m5-1'b1;
												
											end
											end
												else if(display_vga==5'b00101)
										begin
											if(F_pic[m6])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m6<=m6-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m6==0)
												m6<=10'd419;
												else
												m6<=m6-1'b1;
												
											end
											end
												else if(display_vga==5'b00110)
										begin
											if(G_pic[m7])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m7<=m7-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m7==0)
												m7<=10'd419;
												else
												m7<=m7-1'b1;
												
											end
											end
												else if(display_vga==5'b00111)
										begin
											if(H_pic[m8])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m8<=m8-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m8==0)
												m8<=10'd419;
												else
												m8<=m8-1'b1;
												
											end
											end
												else if(display_vga==5'b01000)
										begin
											if(I_pic[m9])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m9<=m9-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m9==0)
												m9<=10'd419;
												else
												m9<=m9-1'b1;
												
											end
											end
												else if(display_vga==5'b01001)
										begin
											if(J_pic[m10])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m10<=m10-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m1==0)
												m10<=10'd419;
												else
												m10<=m10-1'b1;
												
											end
											end
												else if(display_vga==5'b01010)
										begin
											if(K_pic[m11])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m11<=m11-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m11==0)
												m11<=10'd419;
												else
												m11<=m11-1'b1;
												
											end
											end
												else if(display_vga==5'b01011)
										begin
											if(L_pic[m12])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m12<=m12-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m12==0)
												m12<=10'd419;
												else
												m12<=m12-1'b1;
												
											end
											end
												else if(display_vga==5'b01100)
										begin
											if(M_pic[m13])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m13<=m13-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m13==0)
												m13<=10'd419;
												else
												m13<=m13-1'b1;
												
											end
											end
												else if(display_vga==5'b01101)
										begin
											if(N_pic[m14])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m14<=m14-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m14==0)
												m14<=10'd419;
												else
												m14<=m14-1'b1;
												
											end
											end
												else if(display_vga==5'b01110)
										begin
											if(o_pic[m15])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m15<=m15-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m15==0)
												m15<=10'd419;
												else
												m15<=m15-1'b1;
												
											end
											end
												else if(display_vga==5'b10000)
										begin
											if(Q_pic[m16])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m16<=m16-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m16==0)
												m16<=10'd419;
												else
												m16<=m16-1'b1;
												
											end
											end
												else if(display_vga==5'b10001)
										begin
											if(R_pic[m17])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m17<=m17-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m17==0)
												m17<=10'd419;
												else
												m17<=m17-1'b1;
												
											end
											end
												else if(display_vga==5'b10010)
										begin
											if(S_pic[m18])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m18<=m18-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m18==0)
												m18<=10'd419;
												else
												m18<=m18-1'b1;
												
											end
											end
												else if(display_vga==5'b10011)
										begin
											if(T_pic[m19])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd255;
												vga_green<= 8'd25;
												m19<=m19-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m19==0)
												m19<=10'd419;
												else
												m19<=m19-1'b1;
												
											end
											end
												else if(display_vga==5'b10100)
										begin
											if(U_pic[m20])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd255;
												vga_green<= 8'd25;
												m20<=m20-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m20==0)
												m20<=10'd419;
												else
												m20<=m20-1'b1;
												
											end
											end
												else if(display_vga==5'b10101)
										begin
											if(V_pic[m21])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd255;
												m21<=m21-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m21==0)
												m21<=10'd419;
												else
												m21<=m21-1'b1;
												
											end
											end
												else if(display_vga==5'b10110)
										begin
											if(W_pic[m22])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd255;
												m22<=m22-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m22==0)
												m22<=10'd419;
												else
												m22<=m22-1'b1;
												
											end
											end
												else if(display_vga==5'b10111)
										begin
											if(x_pic[m23])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd255;
												m23<=m23-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m23==0)
												m23<=10'd419;
												else
												m23<=m23-1'b1;
												
											end
											end
												else if(display_vga==5'b11000)
										begin
											if(Y_pic[m24])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd255;
												m24<=m24-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m24==0)
												m1<=10'd419;
												else
												m24<=m24-1'b1;
												
											end
											end
												else if(display_vga==5'b11001)
										begin
											if(Z_pic[m25])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd225;
												vga_green<= 8'd25;
												m25<=m25-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m25==0)
												m25<=10'd419;
												else
												m25<=m25-1'b1;
												
											end
											end
												else if(display_vga==5'b01111)
										begin
											if(P_pic[m26])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m26<=m26-1'b1;
											end
											else
											begin
												vga_red<= 8'd0;
												vga_blue<= 8'd0;
												vga_green<= 8'd0;
												if(m26==0)
												m26<=10'd419;
												else
												m26<=m26-1'b1;
												
											end
											end

				else begin
				vga_red<= 8'd127;
				vga_blue<= 8'd158;
				vga_green<= 8'd136;
				end
			end
			else
			begin
				vga_red<= 8'd255;
				vga_blue<= 8'd255;
				vga_green<= 8'd255;				
			end

				if(onn==1'b1)
				begin
					
					//if((pixel_counter >= 10'd0 && pixel_counter <= 10'd210)  && (line_counter >= 10'd0 && line_counter <= 10'd157)) 
					begin
						if((pixel_counter > 10'd30 && pixel_counter <= 10'd60)  && (line_counter > 10'd20 && line_counter <= 10'd34))
						begin
							if(display_vga==5'b00000)
									begin
										vga_red<= 8'd255;
										vga_blue<= 8'd255;
										vga_green<= 8'd255;
										m11<=419;
									end
			
									else if(display_vga==5'b00001)
										begin
											if(A_pic[m1])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m1<=m1-1'b1;
											end
										end
									else if(display_vga==5'b00010)
										begin
											if(B_pic[m2])
											begin
												vga_red<= 8'd255;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m2<=m2-1'b1;
											end
										end	
									else if(display_vga==5'b00011)
										begin
											if(C_pic[m3])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m3<=m3-1'b1;
											end
										end
									else if(display_vga==5'b00100)
										begin
											if(D_pic[m4])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m4<=m4-1'b1;
											end
										end
									else if(display_vga==5'b00101)
										begin
											if(E_pic[m5])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m5<=m5-1'b1;
											end
										end
									else if(display_vga==5'b00110)
										begin
											if(F_pic[m6])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m6<=m6-1'b1;
											end
										end
									else if(display_vga==5'b00111)
										begin
											if(G_pic[m7])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m7<=m7-1'b1;
											end
										end
									else if(display_vga==5'b01000)
										begin
											if(H_pic[m8])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m8<=m8-1'b1;
											end
										end
									else if(display_vga==5'b01001)
										begin
											if(I_pic[m9])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m9<=m9-1'b1;
											end
										end
									else if(display_vga==5'b01010)
										begin
											if(J_pic[m10])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m10<=m10-1'b1;
											end
										end
									else if(display_vga==5'b01011)
										begin
											if(K_pic[m11])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m11<=m11-1'b1;
											end
										end
									else if(display_vga==5'b01100)
										begin
											if(L_pic[m12])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m12<=m12-1'b1;
											end
										end
									else if(display_vga==5'b01101)
										begin
											if(M_pic[m13])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m13<=m13-1'b1;
											end
										end
									else if(display_vga==5'b01110)
										begin
											if(N_pic[m14])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m14<=m14-1'b1;
											end
										end
									else if(display_vga==5'b01111)
										begin
											if(o_pic[m15])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m15<=m15-1'b1;
											end
										end
									else if(display_vga==5'b10000)
										begin
											if(P_pic[m16])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m16<=m16-1'b1;
											end
										end
									else if(display_vga==5'b10001)
										begin
											if(Q_pic[m17])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m17<=m17-1'b1;
											end
										end
									else if(display_vga==5'b10010)
										begin
											if(R_pic[m18])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m18<=m18-1'b1;
											end
										end
									else if(display_vga==5'b10011)
										begin
											if(S_pic[m19])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m19<=m19-1'b1;
											end
										end
									else if(display_vga==5'b10100)
										begin
											if(T_pic[m20])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m20<=m20-1'b1;
											end
										end
									else if(display_vga==5'b10101)
										begin
											if(U_pic[m21])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m21<=m21-1'b1;
											end
										end
									else if(display_vga==5'b10110)
										begin
											if(V_pic[m11])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m22<=m22-1'b1;
											end
										end
									else if(display_vga==5'b10111)
										begin
											if(W_pic[m23])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m23<=m23-1'b1;
											end
										end
									else if(display_vga==5'b11000)
										begin
											if(x_pic[m24])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m24<=m24-1'b1;
											end
										end
									else if(display_vga==5'b11001)
										begin
											if(Y_pic[m25])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m25<=m25-1'b1;
											end
										end
									else if(display_vga==5'b11010)
										begin
											if(Z_pic[m26])
											begin
												vga_red<= 8'd25;
												vga_blue<= 8'd25;
												vga_green<= 8'd25;
												m26<=m26-1'b1;
											end
										end
									
					end
				end
	end	
            /*else
				begin
							vga_red<= 8'd0;
							vga_blue<= 8'd0;
							vga_green<= 8'd255;					
				end*/
	
	end
	end
end
	///////////////////////////////////////////////////////////////////////////////
//Horizontal and Vertical counters

always @ (posedge divcntr)
begin
	if (reset)
	begin
		pixel_counter	<= H_TOTAL - 20; 
		line_counter	<= V_TOTAL - 1; 
	end
	else
	begin
		// last pixel in the line
		if (pixel_counter == (H_TOTAL - 1))
		begin
			pixel_counter <= {PW{1'b0}};
			
			// last pixel in last line of frame
			if (line_counter == (V_TOTAL - 1))
				line_counter <= {LW{1'b0}};
			// last pixel but not last line
			else
				line_counter <= line_counter + LINE_COUNTER_INCREMENT;
		end
		else 
			pixel_counter <= pixel_counter + PIXEL_COUNTER_INCREMENT;  
	end
	
end
///////////////////////////////////////////////////////////////////////////////////////////////////
//End of frame and end of active frame
always @ (posedge divcntr) 
begin
	if (reset)
	begin
		end_of_active_frame <= 1'b0;
		end_of_frame		<= 1'b0;
	end
	else
	begin
		if ((line_counter == (V_ACTIVE - 1)) &&
			(pixel_counter == (H_ACTIVE - 2)))
			end_of_active_frame <= 1'b1;
		else
			end_of_active_frame <= 1'b0;

		if ((line_counter == (V_TOTAL - 1)) && 
			(pixel_counter == (H_TOTAL - 2)))
			end_of_frame <= 1'b1;
		else
			end_of_frame <= 1'b0;
	end
end
		

///////////////////////////////////////////////////////////////////////////////////////////////////
//Sync pulses

always @ (posedge divcntr) 
begin
	if (reset)
	begin
		early_hsync_pulse <= 1'b0;
		early_vsync_pulse <= 1'b0;
		
		hsync_pulse <= 1'b0;
		vsync_pulse <= 1'b0;
		
		csync_pulse	<= 1'b0;
	end
	else
	begin
		// start of horizontal sync
		if (pixel_counter == (H_ACTIVE + H_FRONT_PORCH - 2))
			early_hsync_pulse <= 1'b1;	
		// end of horizontal sync
		else if (pixel_counter == (H_TOTAL - H_BACK_PORCH - 2))
			early_hsync_pulse <= 1'b0;	
			
		// start of vertical sync
		if ((line_counter == (V_ACTIVE + V_FRONT_PORCH - 1)) && 
				(pixel_counter == (H_TOTAL - 2)))
			early_vsync_pulse <= 1'b1;
		// end of vertical sync
		else if ((line_counter == (V_TOTAL - V_BACK_PORCH - 1)) && 
				(pixel_counter == (H_TOTAL - 2)))
			early_vsync_pulse <= 1'b0;
			
		hsync_pulse <= early_hsync_pulse;
		vsync_pulse <= early_vsync_pulse;

		csync_pulse <= early_hsync_pulse ^ early_vsync_pulse;
	end
end


///////////////////////////////////////////////////////////////////////////////////////////////////

// Blanking pulse signals

always @ (posedge divcntr) 
begin
	if (reset)
	begin
		hblanking_pulse	<= 1'b1;
		vblanking_pulse	<= 1'b1;
		
		blanking_pulse	<= 1'b1;
	end
	else
	begin
		if (pixel_counter == (H_ACTIVE - 2))
			hblanking_pulse<= 1'b1;
		else if (pixel_counter == (H_TOTAL - 2))
			hblanking_pulse<= 1'b0;
		
		if ((line_counter == (V_ACTIVE - 1)) &&
				(pixel_counter == (H_TOTAL - 2))) 
			vblanking_pulse<= 1'b1;
		else if ((line_counter == (V_TOTAL - 1)) &&
				(pixel_counter == (H_TOTAL - 2))) 
			vblanking_pulse<= 1'b0;
			
		blanking_pulse<= hblanking_pulse | vblanking_pulse;
	end
end

endmodule
